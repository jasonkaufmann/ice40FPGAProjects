module display (
    input [7:0] data
);

//instantiate a memory block so 
endmodule 